module ChipInterface

(input logic [17:0] SW,
output logic [17:0] LEDR,
output logic [7:0] LEDG,
output logic [6:0] HEX7, HEX6, HEX5, HEX4,
HEX3, HEX2, HEX1, HEX0);
  
//not done
